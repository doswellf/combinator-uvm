//This is dummy DUT. 

module dut_dummy( input apb_clock, input apb_reset, apb_if apb_if);

endmodule
