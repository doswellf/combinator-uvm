//This is dummy DUT. 

module dut_dummy( input clock, input reset, uart_if uart_if0);


endmodule

 
