`ifndef AHB_DEFINES
    `define AHB_DEFINES

    `ifndef AHB_DATA_WIDTH
        `define AHB_DATA_WIDTH 32 // AHB data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH
        `define AHB_ADDR_WIDTH 32 // AHB address bus max width
    `endif
`endif
