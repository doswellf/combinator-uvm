/*-------------------------------------------------------------------------
File name   : spi_defines.svh
Title       : APB - SPI defines
Project     :
Created     :
Description : defines for the APB-SPI Environment
Notes       : 
----------------------------------------------------------------------*/
//   Copyright 1999-2010 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH
`define APB_SPI_DEFINES_SVH

`define SPI_RX0_REG    32'h00
`define SPI_RX1_REG    32'h04
`define SPI_RX2_REG    32'h08
`define SPI_RX3_REG    32'h0C
`define SPI_TX0_REG    32'h00
`define SPI_TX1_REG    32'h04
`define SPI_TX2_REG    32'h08
`define SPI_TX3_REG    32'h0C
`define SPI_CTRL_REG   32'h10
`define SPI_DIV_REG    32'h14
`define SPI_SS_REG     32'h18

`endif
