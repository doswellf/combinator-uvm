/*******************************************************************************
  FILE : apb_types.sv
*******************************************************************************/
//   Copyright 1999-2010 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------


`ifndef APB_TYPES_SVH
`define APB_TYPES_SVH

//------------------------------------------------------------------------------
// apb transfer enums, parameters, and events
typedef enum { APB_READ = 0, APB_WRITE = 1 } apb_direction_enum;

`endif  // APB_TYPES_SVH
